/********************************************************************************
// @project       Object Detection & Tracking Uint(ODTU)
// @filename      sync_bram_sdp.v
// @author        3book
// @description   
// @created       2020-02-10T03:24:19.113Z+08:00
// @copyright     Copyright (c) 2019 
// @last-modified 2020-03-31T22:20:11.792Z+08:00
*******************************************************************************/

`timescale 1ns/100ps
module sync_bram_sdp #(
parameter   WIDTH =144    ,//
parameter   DEPTH =8192,//
parameter   BRAM_SIZE   ="18Kb"      , // Target BRAM, "18Kb" or "36Kb" 
parameter   DEVICE      ="7SERIES"   , // Target device: "7SERIES" 
parameter   DO_REG      =0           ,// Optional output register (0 or 1)
parameter   INIT_FILE   ="NONE"      ,
parameter   SIM_COLLISION_CHECK ="ALL" , // Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
parameter   SRVAL   =72'h000000000000000000, // Set/Reset value for port output
parameter   INIT    =72'h000000000000000000,  // Initial values on output port
parameter   WRITE_MODE  ="WRITE_FIRST"  // Specify "READ_FIRST" for same clock or synchronous clocks
)(
input               clk,// 1-bit input clock
input               rst,// 1-bit input reset
output  [WIDTH-1:0] rddata,// Output read data port, width defined by READ_WIDTH parameter
input   [$clog2(DEPTH)-1:0] rdaddr, // Input read address, width defined by read port depth
input               rden,// 1-bit input read port enable
// input               regce,// 1-bit input read output register enable
input               wren,// 1-bit input write port enable
input   [$clog2(DEPTH)-1:0] wraddr,// Input write address, width defined by write port depth
input   [WIDTH-1:0] wrdata// Input write data port, width defined by WRITE_WIDTH parameter
);

// `define macro_name (arguments) text_string (arguments)
   ///////////////////////////////////////////////////////////////////////
   //  READ_WIDTH | BRAM_SIZE | READ Depth  | RDADDR Width |            //
   // WRITE_WIDTH |           | WRITE Depth | WRADDR Width |  WE Width  //
   // ============|===========|=============|==============|============//
   //    37-72    |  "36Kb"   |      512    |     9-bit    |    8-bit   //
   //    19-36    |  "36Kb"   |     1024    |    10-bit    |    4-bit   //
   //    19-36    |  "18Kb"   |      512    |     9-bit    |    4-bit   //
   //    10-18    |  "36Kb"   |     2048    |    11-bit    |    2-bit   //
   //    10-18    |  "18Kb"   |     1024    |    10-bit    |    2-bit   //
   //     5-9     |  "36Kb"   |     4096    |    12-bit    |    1-bit   //
   //     5-9     |  "18Kb"   |     2048    |    11-bit    |    1-bit   //
   //     3-4     |  "36Kb"   |     8192    |    13-bit    |    1-bit   //
   //     3-4     |  "18Kb"   |     4096    |    12-bit    |    1-bit   //
   //       2     |  "36Kb"   |    16384    |    14-bit    |    1-bit   //
   //       2     |  "18Kb"   |     8192    |    13-bit    |    1-bit   //
   //       1     |  "36Kb"   |    32768    |    15-bit    |    1-bit   //
   //       1     |  "18Kb"   |    16384    |    14-bit    |    1-bit   //
   ///////////////////////////////////////////////////////////////////////
localparam W0 = (BRAM_SIZE=="18Kb") ? 36:72, H0 = 512    ;
localparam W1 = (BRAM_SIZE=="18Kb") ? 18:36, H1 = 1024   ;
localparam W2 = (BRAM_SIZE=="18Kb") ?  9:18, H2 = 2048   ;
localparam W3 = (BRAM_SIZE=="18Kb") ?  4: 9, H3 = 4096   ;
localparam W4 = (BRAM_SIZE=="18Kb") ?  2: 4, H4 = 8192   ;
localparam W5 = (BRAM_SIZE=="18Kb") ?  1: 2, H5 = 16384  ;
localparam W6 = (BRAM_SIZE=="18Kb") ?  1: 1, H6 = (BRAM_SIZE=="18Kb") ? 16384:32768  ;
localparam WN0 = WIDTH/W0 + (WIDTH%W0>0), HN0 = DEPTH/H0 + (DEPTH%H0>0);
localparam WN1 = WIDTH/W1 + (WIDTH%W1>0), HN1 = DEPTH/H1 + (DEPTH%H1>0);
localparam WN2 = WIDTH/W2 + (WIDTH%W2>0), HN2 = DEPTH/H2 + (DEPTH%H2>0);
localparam WN3 = WIDTH/W3 + (WIDTH%W3>0), HN3 = DEPTH/H3 + (DEPTH%H3>0);
localparam WN4 = WIDTH/W4 + (WIDTH%W4>0), HN4 = DEPTH/H4 + (DEPTH%H4>0);
localparam WN5 = WIDTH/W5 + (WIDTH%W5>0), HN5 = DEPTH/H5 + (DEPTH%H5>0);
localparam WN6 = WIDTH/W6 + (WIDTH%W6>0), HN6 = DEPTH/H6 + (DEPTH%H6>0);
localparam N0= WN0*HN0;
localparam N1= WN1*HN1;
localparam N2= WN2*HN2;
localparam N3= WN3*HN3;
localparam N4= WN4*HN4;
localparam N5= WN5*HN5;
localparam N6= WN6*HN6;
localparam RW = N0<N1 ? W0:
                N1<N2 ? W1:
                N2<N3 ? W2:
                N3<N4 ? W3:
                N4<N5 ? W4:
                N5<N6 ? W5:
                        W6;
localparam RH = N0<N1 ? H0:
                N1<N2 ? H1:
                N2<N3 ? H2:
                N3<N4 ? H3:
                N4<N5 ? H4:
                N5<N6 ? H5:
                        H6;
localparam WN = WIDTH/RW + (WIDTH%RW>0);                    
localparam HN = DEPTH/RH + (DEPTH%RH>0);                    
wire [RW*WN-1:0] DI;
wire [RW*WN-1:0] DO;
wire [HN-1:0] ren;
wire [HN-1:0] wen;
wire [$clog2(RH)-1:0] raddr;
wire [$clog2(RH)-1:0] waddr;
assign DI = {{RW*WN-WIDTH{1'b0}},wrdata};
assign rddata = DO[0+:WIDTH];
genvar i,j;
generate 
    if (DEPTH>RH) begin
        assign raddr = rdaddr[0+:$clog2(RH)];
        assign waddr = wraddr[0+:$clog2(RH)];
    end else begin
        assign raddr = rdaddr;
        assign waddr = wraddr;
        // assign raddr = {'b0,rdaddr};
        // assign waddr = {'b0,wraddr};
    end

    for (j=0;j<HN;j=j+1) begin
        localparam [$clog2(HN)-1:1] ADDR_H = j;
        if (DEPTH>RH) begin
            assign ren[j]= (rdaddr[$clog2(DEPTH)-1:$clog2(RH)]==ADDR_H)? rden:1'b0;
            assign wen[j]= (wraddr[$clog2(DEPTH)-1:$clog2(RH)]==ADDR_H)? wren:1'b0;
        end else begin
            assign ren[j]= rden;
            assign wen[j]= wren;
        end
    end
    for (i=0;i<WN;i=i+1) begin:HORIZONTAL
        for (j=0;j<HN;j=j+1) begin:VERTICAL
   BRAM_SDP_MACRO #(
      .BRAM_SIZE(BRAM_SIZE), // Target BRAM, "18Kb" or "36Kb" 
      .DEVICE("7SERIES"), // Target device: "7SERIES" 
      .WRITE_WIDTH(RW),    // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
      .READ_WIDTH(RW),     // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
      .DO_REG(0),         // Optional output register (0 or 1)
      .INIT_FILE ("NONE"),
      .SIM_COLLISION_CHECK ("ALL"), // Collision check enable "ALL", "WARNING_ONLY",
                                    //   "GENERATE_X_ONLY" or "NONE" 
      .SRVAL(72'h000000000000000000), // Set/Reset value for port output
      .INIT(72'h000000000000000000),  // Initial values on output port
      .WRITE_MODE("WRITE_FIRST"),  // Specify "READ_FIRST" for same clock or synchronous clocks
                                   //   Specify "WRITE_FIRST for asynchronous clocks on ports
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),

      // The next set of INIT_xx are valid when configured as 36Kb
      .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),

      // The next set of INITP_xx are for the parity bits
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),

      // The next set of INITP_xx are valid when configured as 36Kb
      .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) BRAM_SDP_MACRO_inst (
      .DO       (DO[i*RW+:RW]           ), // Output read data port, width defined by READ_WIDTH parameter
      .DI       (DI[i*RW+:RW]           ), // Input write data port, width defined by WRITE_WIDTH parameter
      .RDADDR   (raddr  ), // Input read address, width defined by read port depth
      .WRADDR   (waddr  ), // Input write address, width defined by write port depth
      .RDCLK    (clk                    ), // 1-bit input read clock
      .RDEN     (ren[j]                ), // 1-bit input read port enable
      .REGCE    (1'b1                   ), // 1-bit input read output register enable
      .RST      (rst                    ), // 1-bit input reset
      .WE       ({((RW+9-1)/9){1'b1}}     ), // Input write enable, width defined by write port depth
    //   .WE       ({$clog2(RW){1'b1}}     ), // Input write enable, width defined by write port depth
      .WRCLK    (clk                    ), // 1-bit input write clock
      .WREN     (wen[j]                )  // 1-bit input write port enable
   );
   // End of BRAM_SDP_MACRO_inst instantiation
        end
    end
endgenerate
endmodule
